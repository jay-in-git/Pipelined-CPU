module AND(
    input Src1_i,
    input Src2_i,
    output Result_o
);

assign Result_o = Src1_i & Src2_i;

endmodule